module MIPS();

endmodule